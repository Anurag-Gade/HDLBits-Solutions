module top_module (
    input [4:0] a, b, c, d, e, f,
    output [7:0] w, x, y, z );//

    wire [31:0] conc_input;
    assign conc_input = {a, b, c, d, e, f, 2'b11};
    
    assign w = conc_input[31:24];
    assign x = conc_input[23:16];
    assign y = conc_input[15:8];
    assign z = conc_input[7:0];

endmodule
